packageMemory_simu.vhd